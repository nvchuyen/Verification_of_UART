

class base_test extends uvm_test  /* base class*/;
	`uvm_component_utils(base_test);
	
	
endclass : base_test