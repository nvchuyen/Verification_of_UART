//--------------------------------------------
//
//
//
//--------------------------------------------
//
// Class Description
//

package test_lib_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
	
	import env_pkg::*;
	import agent_pkg::*;
	import seq_lib_pkg::*;
	

 // Includes:
`include "base_test.svh"
`include "first_test.svh"
`include "test_rb6l.svh"
`include "test_rb5l.svh"
`include "test_rb7l.svh"
`include "test_rb8l.svh"
`include "test_rb5lwop.svh"
`include "test_rb6lwop.svh"
`include "test_rb7lwop.svh"
`include "test_rb8lwop.svh"

endpackage : test_lib_pkg

